* Netlist before simplification

* cell NET_VSS$2
.SUBCKT NET_VSS$2
.ENDS NET_VSS$2

* cell NET_ENABLE$3
.SUBCKT NET_ENABLE$3
.ENDS NET_ENABLE$3

* cell NET_OUT$3
.SUBCKT NET_OUT$3
.ENDS NET_OUT$3

* cell NET_VDD$3
.SUBCKT NET_VDD$3
.ENDS NET_VDD$3

* cell NET_FB$3
.SUBCKT NET_FB$3
.ENDS NET_FB$3

* cell NET_$10$3
.SUBCKT NET_$10$3
.ENDS NET_$10$3

* cell NET_$9$3
.SUBCKT NET_$9$3
.ENDS NET_$9$3

* cell NET_$8$3
.SUBCKT NET_$8$3
.ENDS NET_$8$3

* cell NET_$7$3
.SUBCKT NET_$7$3
.ENDS NET_$7$3

* cell NET_$6$3
.SUBCKT NET_$6$3
.ENDS NET_$6$3

* cell NET_$5$3
.SUBCKT NET_$5$3
.ENDS NET_$5$3

* cell NET_$4$3
.SUBCKT NET_$4$3
.ENDS NET_$4$3

* cell NET_$3$3
.SUBCKT NET_$3$3
.ENDS NET_$3$3

* cell NET_$2$3
.SUBCKT NET_$2$3
.ENDS NET_$2$3

* cell NET_$1$3
.SUBCKT NET_$1$3
.ENDS NET_$1$3

* cell NET_VSS$1
.SUBCKT NET_VSS$1
.ENDS NET_VSS$1

* cell NET_ENABLE$2
.SUBCKT NET_ENABLE$2
.ENDS NET_ENABLE$2

* cell NET_OUT$2
.SUBCKT NET_OUT$2
.ENDS NET_OUT$2

* cell NET_VDD$2
.SUBCKT NET_VDD$2
.ENDS NET_VDD$2

* cell NET_FB$2
.SUBCKT NET_FB$2
.ENDS NET_FB$2

* cell NET_$10$2
.SUBCKT NET_$10$2
.ENDS NET_$10$2

* cell NET_$9$2
.SUBCKT NET_$9$2
.ENDS NET_$9$2

* cell NET_$8$2
.SUBCKT NET_$8$2
.ENDS NET_$8$2

* cell NET_$7$2
.SUBCKT NET_$7$2
.ENDS NET_$7$2

* cell NET_$6$2
.SUBCKT NET_$6$2
.ENDS NET_$6$2

* cell NET_$5$2
.SUBCKT NET_$5$2
.ENDS NET_$5$2

* cell NET_$4$2
.SUBCKT NET_$4$2
.ENDS NET_$4$2

* cell NET_$3$2
.SUBCKT NET_$3$2
.ENDS NET_$3$2

* cell NET_$2$2
.SUBCKT NET_$2$2
.ENDS NET_$2$2

* cell NET_$1$2
.SUBCKT NET_$1$2
.ENDS NET_$1$2

* cell NET_VSS
.SUBCKT NET_VSS
.ENDS NET_VSS

* cell NET_ENABLE$1
.SUBCKT NET_ENABLE$1
.ENDS NET_ENABLE$1

* cell NET_OUT$1
.SUBCKT NET_OUT$1
.ENDS NET_OUT$1

* cell NET_VDD$1
.SUBCKT NET_VDD$1
.ENDS NET_VDD$1

* cell NET_FB$1
.SUBCKT NET_FB$1
.ENDS NET_FB$1

* cell NET_$10$1
.SUBCKT NET_$10$1
.ENDS NET_$10$1

* cell NET_$9$1
.SUBCKT NET_$9$1
.ENDS NET_$9$1

* cell NET_$8$1
.SUBCKT NET_$8$1
.ENDS NET_$8$1

* cell NET_$7$1
.SUBCKT NET_$7$1
.ENDS NET_$7$1

* cell NET_$6$1
.SUBCKT NET_$6$1
.ENDS NET_$6$1

* cell NET_$5$1
.SUBCKT NET_$5$1
.ENDS NET_$5$1

* cell NET_$4$1
.SUBCKT NET_$4$1
.ENDS NET_$4$1

* cell NET_$3$1
.SUBCKT NET_$3$1
.ENDS NET_$3$1

* cell NET_$2$1
.SUBCKT NET_$2$1
.ENDS NET_$2$1

* cell NET_$1$1
.SUBCKT NET_$1$1
.ENDS NET_$1$1

* cell NET_BULK,VSS
.SUBCKT NET_BULK,VSS
.ENDS NET_BULK,VSS

* cell NET_VDD
.SUBCKT NET_VDD
.ENDS NET_VDD

* cell NET_$2
.SUBCKT NET_$2
.ENDS NET_$2

* cell NET_ENABLE
.SUBCKT NET_ENABLE
.ENDS NET_ENABLE

* cell NET_OUT
.SUBCKT NET_OUT
.ENDS NET_OUT

* cell NET_FB
.SUBCKT NET_FB
.ENDS NET_FB

* cell NET_$10
.SUBCKT NET_$10
.ENDS NET_$10

* cell NET_$9
.SUBCKT NET_$9
.ENDS NET_$9

* cell NET_$8
.SUBCKT NET_$8
.ENDS NET_$8

* cell NET_$7
.SUBCKT NET_$7
.ENDS NET_$7

* cell NET_$6
.SUBCKT NET_$6
.ENDS NET_$6

* cell NET_$5
.SUBCKT NET_$5
.ENDS NET_$5

* cell NET_$4
.SUBCKT NET_$4
.ENDS NET_$4

* cell NET_$3
.SUBCKT NET_$3
.ENDS NET_$3

* cell NET_$1
.SUBCKT NET_$1
.ENDS NET_$1

* cell NET_$I3$3
.SUBCKT NET_$I3$3
.ENDS NET_$I3$3

* cell NET_$I3$2
.SUBCKT NET_$I3$2
.ENDS NET_$I3$2

* cell NET_$I3$1
.SUBCKT NET_$I3$1
.ENDS NET_$I3$1

* cell NET_$I3
.SUBCKT NET_$I3
.ENDS NET_$I3

* cell RINGO
.SUBCKT RINGO
* net 11 FB
* net 12 VDD
* net 13 OUT
* net 14 ENABLE
* net 15 VSS
* cell instance $1 r0 *1 1.8,0
X$1 12 1 15 12 11 14 15 ND2X1
* cell instance $2 r0 *1 4.2,0
X$2 12 2 15 12 1 15 INVX1
* cell instance $3 r0 *1 6,0
X$3 12 3 15 12 2 15 INVX1
* cell instance $4 r0 *1 7.8,0
X$4 12 4 15 12 3 15 INVX1
* cell instance $5 r0 *1 9.6,0
X$5 12 5 15 12 4 15 INVX1
* cell instance $6 r0 *1 11.4,0
X$6 12 6 15 12 5 15 INVX1
* cell instance $7 r0 *1 13.2,0
X$7 12 7 15 12 6 15 INVX1
* cell instance $8 r0 *1 15,0
X$8 12 8 15 12 7 15 INVX1
* cell instance $9 r0 *1 16.8,0
X$9 12 9 15 12 8 15 INVX1
* cell instance $10 r0 *1 18.6,0
X$10 12 10 15 12 9 15 INVX1
* cell instance $11 r0 *1 20.4,0
X$11 12 11 15 12 10 15 INVX1
* cell instance $12 r0 *1 22.2,0
X$12 12 13 15 12 11 15 INVX1
* cell instance $13 r0 *1 3.28,4
X$13 11 M1M2
* cell instance $14 r0 *1 21.42,4
X$14 11 M1M2
* cell instance $15 r0 *1 0.6,0
X$15 12 15 TIE
* cell instance $16 r0 *1 0,0
X$16 12 15 12 EMPTY
* cell instance $17 r0 *1 24,0
X$17 12 15 TIE
* cell instance $18 r0 *1 25.2,0
X$18 12 15 12 EMPTY
* cell instance $19 r0 *1 23.6,4
X$19 13 M1M2
* cell instance $20 r0 *1 2.6,3.1
X$20 14 M1M2
.ENDS RINGO

* cell INVX1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin IN
* pin BULK
.SUBCKT INVX1 1 2 3 4 5 6
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 IN
* net 6 BULK
* cell instance $1 r0 *1 0.3,5.05
X$1 5 2 1 PMOS3
* cell instance $2 r0 *1 0.3,1.66
X$2 5 2 3 NMOS2
* cell instance $3 r0 *1 0.6,3.1
X$3 5 POLYM1
* device instance $1 r0 *1 0.85,5.8 LVPMOS
M$1 1 5 2 4 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.6375P PS=3.85U PD=3.85U
* device instance $2 r0 *1 0.85,2.135 LVNMOS
M$2 3 5 2 6 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.40375P PS=2.75U PD=2.75U
.ENDS INVX1

* cell EMPTY
* pin 
* pin 
* pin 
.SUBCKT EMPTY 1 2 3
.ENDS EMPTY

* cell TIE
* pin VDD
* pin VSS
.SUBCKT TIE 1 2
* net 1 VDD
* net 2 VSS
.ENDS TIE

* cell M1M2
* pin 
.SUBCKT M1M2 1
.ENDS M1M2

* cell ND2X1
* pin VDD
* pin OUT
* pin VSS
* pin 
* pin B
* pin A
* pin BULK
.SUBCKT ND2X1 1 2 3 4 5 6 7
* net 1 VDD
* net 2 OUT
* net 3 VSS
* net 5 B
* net 6 A
* net 7 BULK
* cell instance $1 r0 *1 0.3,5.05
X$1 6 1 2 PMOS3
* cell instance $2 r0 *1 1,5.05
X$2 5 2 1 PMOS3
* cell instance $3 r0 *1 1,1.66
X$3 5 2 8 NMOS2
* cell instance $4 r0 *1 0.3,1.66
X$4 6 8 3 NMOS2
* cell instance $5 r0 *1 1.48,4
X$5 5 POLYM1
* cell instance $6 r0 *1 0.8,3.1
X$6 6 POLYM1
* device instance $1 r0 *1 0.85,5.8 LVPMOS
M$1 2 6 1 4 LVPMOS L=0.25U W=1.5U AS=0.6375P AD=0.3375P PS=3.85U PD=1.95U
* device instance $2 r0 *1 1.55,5.8 LVPMOS
M$2 1 5 2 4 LVPMOS L=0.25U W=1.5U AS=0.3375P AD=0.6375P PS=1.95U PD=3.85U
* device instance $3 r0 *1 0.85,2.135 LVNMOS
M$3 3 6 8 7 LVNMOS L=0.25U W=0.95U AS=0.40375P AD=0.21375P PS=2.75U PD=1.4U
* device instance $4 r0 *1 1.55,2.135 LVNMOS
M$4 8 5 2 7 LVNMOS L=0.25U W=0.95U AS=0.21375P AD=0.40375P PS=1.4U PD=2.75U
.ENDS ND2X1

* cell PMOS3
* pin 
* pin 
* pin 
.SUBCKT PMOS3 1 2 3
.ENDS PMOS3

* cell NMOS2
* pin 
* pin 
* pin 
.SUBCKT NMOS2 1 2 3
.ENDS NMOS2

* cell POLYM1
* pin 
.SUBCKT POLYM1 1
.ENDS POLYM1
